module gnd_circuit(
   output out
);
	assign out = 1'b0;
endmodule 