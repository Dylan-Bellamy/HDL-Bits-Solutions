module wire_circuit(
   input in,
   output out
);
	assign out = in;	
endmodule 