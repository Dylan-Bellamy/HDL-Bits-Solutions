module zero_module ( zero );
	output zero;
	assign zero = 0;
endmodule 